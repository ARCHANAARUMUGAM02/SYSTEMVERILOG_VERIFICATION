interface inter;
  logic clk;
  logic we;
  logic[3:0]addr;
  logic[7:0]din;
  logic[7:0]dout;
endinterface
  
