interface inter();
  bit clk;
  logic rst;
  logic rd_en;
  logic wr_en;
  logic full,empty;
  logic[8:0] din;
  logic[7:0] dout;
endinterface
  
  
